`ifndef DEFINES
`define DEFINES

`endif // DEFINES
