/*
 * Joseph Ravichandran
 * December 6, 2020
 */

/*
 * psp
 * A pretty secure processor.
 */
module psp
    (
        input logic clk
    );

    // Main Memory

    // Caches

    // Core

endmodule
